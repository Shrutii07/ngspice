*bandpassfilter opamp
.include LF356.MOD
V1  1 0     DC 0 AC 1
C1  1 p1    10n
R1  p1 0    7.23431K

R2  n1 0    10K
R3  n1 4    10K

R4  4 p2    2.2105K
C2  p2 0    10n

R5  n2 0    10K
R6  n2 out  10K
RL  out 0   10G

Vcc vp 0    DC 12
Vee vn 0    DC -12

X1  p1 n1 vp vn 4  LF356/NS  
X2  p2 n2 vp vn out LF356/NS

.ac dec 100 1 1Meg   * AC sweep from 100Hz to 1MHz in steps of 1Hz
.control
run
plot db(v(out))
.endc
.end
