D Flip Flop

vclk clk 0 PULSE(0 5 0 0 0 5m 10m)
vd d 0 PULSE(0 9.9 0 0 0 7m 14m)

.subckt not 1 2
	v1 3 0 5
	m1 3 1 2 3 PFET
	m3 2 1 0 0 NFET

	.model PFET PMOS
	.model NFET NMOS
.ends

.subckt flipFlop d clk q notq
	vdd vd 0 5

	Xu1 clk ntclk not

	mp1 vd d n1 vd PFET
	mp2 n1 ntclk notq vd PFET

	mn1 notq clk n2 0 NFET
	mn2 n2 d 0 0 NFET


	mp3 vd notq q vd PFET

	mn3 q notq 0 0 NFET


	mp4 vd q n3 vd PFET
	mp5 n3 clk notq vd PFET

	mn4 notq ntclk n4 0 NFET
	mn5 n4 q 0 0 NFET


	.model PFET PMOS
	.model NFET NMOS
.ends

Xu1 d clk q notq flipFlop

.tran 1u 80m
.control
run

set color0=black
set color1=white
set color2=red
set color3=blue
set color4=green
set color5 = violet

plot v(clk) v(d)+10 v(q)+25 v(notq)+40 

.endc
.end
