*Chua circuit using transistor

l1 1 0 8.5m
c2 1 0 47n
r9 1 2 1.6k
c1 2 0 4.6n

d1 3 2 
r3 3 0 3.3k
r2 3 6 47k
v1 0 6 dc 9v
d2 2 4 
r1 4 0 3.3k
r4 4 7 47k
v2 7 0 dc 9v
r7 2 5 290
r6 5 11 290
q1 8 8 6 bjtn
q2 9 9 7 bjtp
q3 9 2 10 bjtn
q4 5 11 10 bjtn
q5 10 8 6 bjtn
q6 5 9 7 bjtp
r8 7 8 5k
r5 11 0 1.2k

.model bjtn npn
.model bjtp pnp

.tran 1u 100m
.control
SET COLOR0 = white
SET COLOR1 = black
SET COLOR2= red
SET COLOR3= blue
SET COLOR4 = brown
Set XbrushWidth = 2
run
plot v(1) vs v(2)
plot v(1) V(2)
linearize
fft V(1) V(2)
plot V(1) V(2) xlimit 0 20kHz
.endc
.end
