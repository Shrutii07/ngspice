* common gate amplifier MOSFET

Vin 1 0 sine(0 4 350)
*Vin 1 0 dc=0 ac=5
C1 1 s1 100u
Rs s1 0 10K

Vdd 2 0 DC 1V
Rd 2 d1 50k
C2 d1 op 100u
Rl op 0 100k

R1 2 g 100K
R2 g 0 1K
Cg g 0 100u

*MX nd ng ns nb mname
M1 d1 g s1 s1 Mos_Shru
.model Mos_Shru NMOS

.tran 1u 10m
* unmcomment above one for transient analysis
* uncomment below one for ac analysis	
*.ac dec 100 1 1Mega

.control
run

plot v(1) v(op)
* unmcomment above one for ip op plot
* uncomment below one for gain plot	
*plot db(v(op))

.endc
.end
