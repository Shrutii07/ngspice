*low-passfilterr opamp

.include LF356.MOD
vin 1 0 dc 0 ac 1

r1 1 2 10K
c1 2 0 100n
r2 3 0 1K
rf 3 4 9K

vcc 5 0 12
vdd 6 0 -12

XU1 2 3 5 6 4 LF356/NS

.ac dec 100 1 1Meg
.control
run
plot vdb(4) 17 xlog
.endc
.end
