*tflipflop
* xor cmos
.subckt XOR n1 n2 b3
	.model NFET NMOS
	.model PFET PMOS
	m1 d1 n1 b1 d1 PFET
	m2 b1 n1 0 0 NFET
	m3 n1 n2 b3 d1 PFET
	m4 b3 n2 0 0 NFET
.ends

*Edge-trigerred D-Flip flop
	*NAND
	.subckt NAND n1 n2 d1
		Vdc dc 0 10
		m1 d1 n1 s1 0 NFET
		m2 s1 n2 0 0 NFET
		m3 dc n1 d1 dc PFET
		m4 dc n2 d1 dc PFET
		.model NFET NMOS
		.model PFET PMOS
	.ends

	*NAND3IP USING 2IPNAND
	.subckt NAND3 in1 in2 in3 out3
		X1 in1 in2 out1 NAND
		X2 out1 out1 out2 NAND
		X3 in3 out2 out3 NAND
	.ends
	.subckt Dflipflop A C Q Qbar
		X1 p4 p1 p3 NAND
		X2 C p3 p1 NAND
		X3 p1 C p4 p2 NAND3
		X4 p2 A p4 NAND
		X5 p1 Qbar Q NAND
		X6 p2 Q Qbar NAND
	.ends

Va A 0 PULSE(9.9 0 1us 1us 1us 20ms 45ms)
Vcin C 0 PULSE(0 9.9 1us 1us 1us 10ms 20ms)
X1 A Q D XOR
X2 D C Q Qbar Dflipflop
.control
tran 0.01ms 90ms
Set Xbrushwidth=2
plot V(C) V(A)+20 V(Q)+40 V(Qbar)+60
.endc
.end
