*Edge_trigerred D-Flip flop

*NAND
.subckt NAND n1 n2 d1
	Vdc dc 0 10
	m1 d1 n1 s1 0 NFET
	m2 s1 n2 0 0 NFET
	m3 dc n1 d1 dc PFET
	m4 dc n2 d1 dc PFET
	.model NFET NMOS
	.model PFET PMOS
.ends

*NAND3IP USING 2IPNAND
.subckt NAND3 in1 in2 in3 out3
	X1 in1 in2 out1 NAND
	X2 out1 out1 out2 NAND
	X3 in3 out2 out3 NAND
.ends

Va A 0 PULSE(0 9.9 1us 1us 1us 10ms 20ms)
Vcin C 0 PULSE(9.9 0 1us 1us 1us 15ms 45ms)

X1 p4 p1 p3 NAND
X2 C p3 p1 NAND
X3 p1 C p4 p2 NAND3
X4 p2 A p4 NAND
X5 p1 Qbar Q NAND
X6 p2 Q Qbar NAND

.control
tran 0.01ms 90ms
Set Xbrushwidth=2
plot V(C) V(A)+20 V(Q)+40 V(Qbar)+60
.endc
.end
