*divider ckt analysis
R1 1 2 1K 
R2 2 0 2K
vin 1 0 dc 5 
.dc vin 0 5.0 0.25 
.control 
run 
plot v(2)
plot v(1,2) 
plot v(1) 
plot v(2)/1K 
plot v(1,2)/1K 
.endc 
.end
