*fullwave rectifier RC

v1 n1 n2 sin(0 2 100)

D1 n1 3 D_shru
D2 n2 3 D_shru
D3 0 n1 D_shru
D4 0 n2 D_shru
R 3 0 1K
C 3 0 9.9uF

.model D_shru D
.tran 10us 10ms	*step of 10usec, total time of 10msec
.control
run
plot v(3)
plot v(n1,n2)
.options savecurrents
plot @C[i] + @R[i]
.endc
.end
