* Colpritt oscillator at 2.2 kHz
.MODEL NPN_Shru npn is=1e-15

Vb  4 0 DC 9

Q1  1 5 2 NPN_Shru

Rc  1 4    5K
Re  2 0    2.7K
Ce  2 0    10u
Ra  4 5    10K
Rb  5 0    4.7K
Cb  5 7    10u
R2  5 7    1M

Co  1 3  10u
C1  3 0  24n
Lt  3 7  240m
C2  7 0  240n

.tran 1u 5000u 20u *Transient response in steps of 1uS, from 20uS to 5000uS
.control
run		
plot v(3)
.endc		
.end



